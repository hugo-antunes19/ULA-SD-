----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Hugo Antunes, Giovanni e Bernardo Pozzato
-- 
-- Create Date:    31/10/2023
-- Module Name:    countertest - Behavioral 
----------------------------------------------------------------------------------
-- Notas: 
-- Fizemos esse arquivo como teste para simular o clock e o contador corretamente
-- Os testes realizados serão anexados devidamente no relatório.
--------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY counter_test IS
END counter_test;
 
ARCHITECTURE behavior OF counter_test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT counter
    PORT(
         selector : IN  std_logic_vector(2 downto 0);
         clk : IN  std_logic;
         step : OUT  std_logic_vector(1 downto 0);
         leds : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

	--Inputs
	
   signal selector : std_logic_vector(2 downto 0) := (others => '0');
   signal clk : std_logic := '0';

	--Outputs

   signal step : std_logic_vector(1 downto 0);
   signal leds : std_logic_vector(3 downto 0);

   	-- Clock period definitions

   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: counter PORT MAP (
          selector => selector,
          clk => clk,
          step => step,
          leds => leds
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait;
   end process;

END;
